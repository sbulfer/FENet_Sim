../../../FENet_Verilog/Interfaces/macCtrlIntf.sv