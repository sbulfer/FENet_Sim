../../FENet_Verilog/Gray_Counter.sv