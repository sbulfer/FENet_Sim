../../../FENet_Verilog/PortConnections/macPort.sv