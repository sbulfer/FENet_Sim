../../../FENet_Verilog/Interfaces/macIntfAr.sv