../../FENet_Verilog/CLK_domain_interface.sv