../../FENet_Verilog/multBus.sv