../../FENet_Verilog/FENet_Module.sv