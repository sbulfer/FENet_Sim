../../FENet_Verilog/FENet_Master.sv