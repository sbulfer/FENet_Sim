../../FENet_Verilog/multBusDecoder.sv