../../FENet_Verilog/Debug_Port.sv