../../TestBenches/FENet_tb.sv