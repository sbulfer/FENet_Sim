../../FENet_Verilog/FENet_Control.sv