../../../FENet_Verilog/Interfaces/procIntf.sv