../../FENet_Verilog/Data_Interface.sv