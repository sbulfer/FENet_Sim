../../FENet_Verilog/Mac_Clk_Gen.sv