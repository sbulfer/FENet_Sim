../../../FENet_Verilog/Interfaces/macClkGenIntf.sv