../../FENet_Verilog/MAC.sv