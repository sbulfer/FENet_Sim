../../../FENet_Verilog/Interfaces/macMstrCtrlIntf.sv