../../FENet_Verilog/Definitions.sv