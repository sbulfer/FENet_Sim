../../../FENet_Verilog/Interfaces/procCtrlIntf.sv