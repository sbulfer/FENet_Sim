../../FENet_Verilog/Cache_Write_Bus.sv