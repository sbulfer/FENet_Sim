../../../FENet_Verilog/PortConnections/ctrlPort.sv