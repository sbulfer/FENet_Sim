../../FENet_Verilog/Scheduler.sv