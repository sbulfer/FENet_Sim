../../../FENet_Verilog/Interfaces/macIntf.sv