../../FENet_Verilog/SRAM.sv