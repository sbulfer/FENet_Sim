../../FENet_Verilog/FPGA_Wrapper.sv