../../../FENet_Verilog/Interfaces/femIntfAr.sv