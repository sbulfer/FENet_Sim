../../../FENet_Verilog/Interfaces/femIntf.sv