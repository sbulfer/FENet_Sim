../../FENet_Verilog/Feature_Engineering_Module.sv