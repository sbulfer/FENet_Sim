../../FENet_Verilog/Input_Queue.sv