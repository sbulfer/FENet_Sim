../../../FENet_Verilog/PortConnections/memPort.sv