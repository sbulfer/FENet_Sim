../../FENet_Verilog/MAC_ctrl.sv