../../FENet_Verilog/External_Interface.sv